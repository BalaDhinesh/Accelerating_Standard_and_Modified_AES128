module MIX_COLUMNS(
    input clk,
    input [127:0] IN_DATA,
    output [127:0] MIXED_DATA
);

reg [127:0] MIXED_DATA_REG;

  always @(*) begin
    MIXED_DATA_REG[127:120] = MIXCOLUMN(IN_DATA[127:120],IN_DATA[119:112],IN_DATA[111:104],IN_DATA[103:96]);
    MIXED_DATA_REG[119:112] = MIXCOLUMN(IN_DATA[119:112],IN_DATA[111:104],IN_DATA[103:96],IN_DATA[127:120]);
    MIXED_DATA_REG[111:104] = MIXCOLUMN(IN_DATA[111:104],IN_DATA[103:96],IN_DATA[127:120],IN_DATA[119:112]);
    MIXED_DATA_REG[103:96] = MIXCOLUMN(IN_DATA[103:96],IN_DATA[127:120],IN_DATA[119:112],IN_DATA[111:104]);

    MIXED_DATA_REG[95:88] = MIXCOLUMN(IN_DATA[95:88],IN_DATA[87:80],IN_DATA[79:72],IN_DATA[71:64]);
    MIXED_DATA_REG[87:80] = MIXCOLUMN(IN_DATA[87:80],IN_DATA[79:72],IN_DATA[71:64],IN_DATA[95:88]);
    MIXED_DATA_REG[79:72] = MIXCOLUMN(IN_DATA[79:72],IN_DATA[71:64],IN_DATA[95:88],IN_DATA[87:80]);
    MIXED_DATA_REG[71:64] = MIXCOLUMN(IN_DATA[71:64],IN_DATA[95:88],IN_DATA[87:80],IN_DATA[79:72]);

    MIXED_DATA_REG[63:56] = MIXCOLUMN(IN_DATA[63:56],IN_DATA[55:48],IN_DATA[47:40],IN_DATA[39:32]);
    MIXED_DATA_REG[55:48] = MIXCOLUMN(IN_DATA[55:48],IN_DATA[47:40],IN_DATA[39:32],IN_DATA[63:56]);
    MIXED_DATA_REG[47:40] = MIXCOLUMN(IN_DATA[47:40],IN_DATA[39:32],IN_DATA[63:56],IN_DATA[55:48]);
    MIXED_DATA_REG[39:32] = MIXCOLUMN(IN_DATA[39:32],IN_DATA[63:56],IN_DATA[55:48],IN_DATA[47:40]);

    MIXED_DATA_REG[31:24] = MIXCOLUMN(IN_DATA[31:24],IN_DATA[23:16],IN_DATA[15:8],IN_DATA[7:0]);
    MIXED_DATA_REG[23:16] = MIXCOLUMN(IN_DATA[23:16],IN_DATA[15:8],IN_DATA[7:0],IN_DATA[31:24]);
    MIXED_DATA_REG[15:8] = MIXCOLUMN(IN_DATA[15:8],IN_DATA[7:0],IN_DATA[31:24],IN_DATA[23:16]);
    MIXED_DATA_REG[7:0] = MIXCOLUMN(IN_DATA[7:0],IN_DATA[31:24],IN_DATA[23:16],IN_DATA[15:8]);
end

assign MIXED_DATA = MIXED_DATA_REG;
   
function [7:0] MIXCOLUMN;
input [7:0] IN1, IN2, IN3, IN4;
    begin
        MIXCOLUMN[7] = IN1[6]^IN2[6]^IN2[7]^IN3[7]^IN4[7];
        MIXCOLUMN[6] = IN1[5]^IN2[5]^IN2[6]^IN3[6]^IN4[6];
        MIXCOLUMN[5] = IN1[4]^IN2[4]^IN2[5]^IN3[5]^IN4[5];
        MIXCOLUMN[4] = IN1[3]^IN1[7]^IN2[3]^IN2[4]^IN2[7]^IN3[4]^IN4[4];
        MIXCOLUMN[3] = IN1[2]^IN1[7]^IN2[2]^IN2[3]^IN2[7]^IN3[3]^IN4[3];
        MIXCOLUMN[2] = IN1[1]^IN2[1]^IN2[2]^IN3[2]^IN4[2];
        MIXCOLUMN[1] = IN1[0]^IN1[7]^IN2[0]^IN2[1]^IN2[7]^IN3[1]^IN4[1];
        MIXCOLUMN[0] = IN1[7]^IN2[7]^IN2[0]^IN3[0]^IN4[0];
    end
endfunction

endmodule